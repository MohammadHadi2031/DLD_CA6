`timescale 1ns/1ns 

module multiplyer (output [31:0]mul, input[15:0] A, B);
assign mul = A * B;
endmodule
